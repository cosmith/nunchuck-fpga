-- 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity FSMAddressTest is
end FSMAddressTest;

architecture Behavioral of FSMAddressTest is

begin


end Behavioral;
